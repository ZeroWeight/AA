module FCore (clk,in,led,num,dot);
input clk;
input in;
output [2:0] led;
output [3:0] num;
output dot;
always @ (posedge in)
begin
end
endmodule
